library verilog;
use verilog.vl_types.all;
entity single_clk_cnt is
end single_clk_cnt;
